`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:   15:53:54 10/28/2019
// Design Name:   ExtendSign
// Module Name:   E:/3rd year/COA Lab/KGP_RISC/extendSign_tb.v
// Project Name:  KGP_RISC
// Target Device:  
// Tool versions:  
// Description:
//
// Verilog Test Fixture created by ISE for module: ExtendSign
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
////////////////////////////////////////////////////////////////////////////////

module extendSign_tb;

// Inputs
reg [15:0] in;

// Outputs
wire [31:0] out;

// Instantiate the Unit Under Test (UUT)
ExtendSign uut (
.in(in),
.out(out)
);

initial begin
// Initialize Inputs
in = 0;

// Wait 100 ns for global reset to finish
#100;
in=16'b1001000100010001;

       
// Add stimulus here

end
     
endmodule